module CommMaster 
	(TX, cmd, snd_cmd, data, clk, rst_n);

///////////////////////////////////////////////
// Module Interface Input and Outputs /////////
///////////////////////////////////////////////

//outputs
output logic TX;

//inputs 
input clk, rst_n;
input [7:0] cmd;
input snd_cmd;
input [15:0] data;


///////////////////////////////////////////////
/// internal signals                        ///
///////////////////////////////////////////////

logic [1:0] sel;
logic trmt;
logic tx_done;
logic frm_snt;
logic set_cmplt, clr_cmplt;

logic [7:0] tx_data; //input to UART
logic [7:0] low_bits, mid_bits;


//// Define state as enumerated type /////
typedef enum reg {IDLE, WAITH, WAITM, WAITL} state_t;
state_t state, nxt_state;


//// instantiate transceiver ////
UART_tx txmod(
	.clk(clk),
	.rst_n(rst_n),
	.TX(TX),
	.trmt(trmt),
	.tx_data(tx_data),
	.tx_done(tx_done));


//// flops for high and mid bits ////
always_ff @(posedge clk) begin
	if(snd_cmd)
		low_bits <= data[7:0];
end

always_ff @(posedge clk) begin
	if(snd_cmd)
		mid_bits <= data[15:8];
end

//// tx_data select logic /////
assign tx_data = 
(sel ==  2'b01) ? mid_bits : 
(sel ==  2'b10) ? cmd[7:0] :
(sel ==  2'b00) ? low_bits; 

always_comb begin 
	sel = 2'b10;
	trmt = 0;
	set_cmplt = 0;
	clr_cmplt = 0;

	case (state)
		IDLE: begin 
			if(snd_cmd) begin
				trmt = 1;
				clr_cmplt = 1;
				sel = 2'b10;
				nxt_state = WAITH;
			end else begin
				nxt_state = IDLE;
			end
		end

		WAITH: begin
			if(tx_done) begin 
				sel = 2'b01;
				trmt = 1;
				nxt_state = WAITM;
			end else begin 
				nxt_state = WAITH;
				sel = 2'b10;
			end
		end

		WAITM: begin
			if(tx_done) begin
				sel = 2'b00;
				trmt = 1;
				nxt_state = WAITL;
			end else begin
				sel = 2'b01;
				nxt_state = WAITM;
			end

		end

	default : begin //WAITL STATE
		if(tx_done) begin
			set_cmplt = 1;
			nxt_state = IDLE;
		end else begin
			nxt_state = WAITL;
			sel = 2'b00;
		end
	end
endcase

end



////////////////////////////
// Infer state flop next //
//////////////////////////
always_ff @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		state <= IDLE;
	else
	state <= nxt_state;
end

endmodule