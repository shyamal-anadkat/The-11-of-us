module tb_tasks ();

endmodule